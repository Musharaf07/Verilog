//Number Sequence in Diamond Pattern Tb
module seq_shape_tb;
  seq_shape duv();
   initial begin
     $display("Sequence Diamond shape:");
     #100;$finish;
     end
 endmodule
